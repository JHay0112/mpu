-- Logic package
-- Defines key logical components such as control and ALU.
--
-- Author: J. L. Hay


library ieee;
use ieee.std_logic_1164.all;

library work;
use work.config.all;


package logic is 
    
    

end package;
