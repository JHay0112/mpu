-- Logic package
-- Defines key logical components such as control and ALU.
--
-- Author: J. L. Hay

library ieee;
use ieee.std_logic_1164.all;

package memory is 

    -- Control logic configuration
    

    -- Control logic specification
    component control is
    
    end component;
    
    -- ALU configuration
    
    
    -- ALU specification
    component alu is
        
    end component;

end package memory;
