-- Arithmetic Logic Unit
--
-- Author: J. L. Hay

library ieee;
use ieee.std_logic_1164.all;

entity alu is 

end alu;

architecture Behavioral of alu is

begin


end Behavioral;
