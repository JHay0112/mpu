-- Control Logic
-- To be implemented as a finite state machine.
--
-- Author: J. L. Hay

library ieee;
use ieee.std_logic_1164.all;

entity control is

end control;

architecture Behavioral of control is

begin


end Behavioral;
