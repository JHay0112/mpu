-- RISC-V Microprocessor
--
-- Author: J. L. Hay

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.config.all;

entity main is
    
end main;

architecture Structural of main is

  

begin



end Structural;
