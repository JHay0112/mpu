-- Device configuration
-- Defines values that defined key properties of the device
-- i.e. the word width
--
-- Author: J. L. Hay

package config is 

    constant WORD_WIDTH : integer := 16;

end package;